magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< locali >>
rect 1371 3292 2927 3621
<< metal1 >>
rect 1501 4304 2805 5234
rect 1382 3717 2805 4149
rect 1382 3045 1639 3717
rect 1884 3045 2141 3717
rect 2548 3045 2805 3717
rect 2231 2940 2246 3010
rect 0 583 14 705
rect 2104 418 2127 555
use cascode_PMOS  cascode_PMOS_0
timestamp 1634927741
transform 1 0 174 0 1 0
box -174 66 5531 3553
use sky130_fd_pr__res_high_po_0p69_D8BZCP  sky130_fd_pr__res_high_po_0p69_D8BZCP_0
timestamp 1634927741
transform 1 0 2149 0 1 4218
box -804 -657 804 657
<< labels >>
rlabel metal1 s 2239 5234 2239 5234 4 VDD
port 1 nsew
rlabel metal1 s 2115 418 2115 418 4 G1
port 2 nsew
rlabel metal1 s 0 638 0 638 4 G2
port 3 nsew
rlabel metal1 s 2238 3010 2238 3010 4 S1
port 4 nsew
<< end >>
