magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< metal4 >>
rect -3351 2998 3351 3100
rect -3351 2762 3095 2998
rect 3331 2762 3351 2998
rect -3351 2678 3351 2762
rect -3351 2442 3095 2678
rect 3331 2442 3351 2678
rect -3351 2358 3351 2442
rect -3351 2122 3095 2358
rect 3331 2122 3351 2358
rect -3351 2038 3351 2122
rect -3351 1802 3095 2038
rect 3331 1802 3351 2038
rect -3351 1718 3351 1802
rect -3351 1482 3095 1718
rect 3331 1482 3351 1718
rect -3351 1398 3351 1482
rect -3351 1162 3095 1398
rect 3331 1162 3351 1398
rect -3351 1078 3351 1162
rect -3351 842 3095 1078
rect 3331 842 3351 1078
rect -3351 758 3351 842
rect -3351 522 3095 758
rect 3331 522 3351 758
rect -3351 438 3351 522
rect -3351 202 3095 438
rect 3331 202 3351 438
rect -3351 118 3351 202
rect -3351 -118 3095 118
rect 3331 -118 3351 118
rect -3351 -202 3351 -118
rect -3351 -438 3095 -202
rect 3331 -438 3351 -202
rect -3351 -522 3351 -438
rect -3351 -758 3095 -522
rect 3331 -758 3351 -522
rect -3351 -842 3351 -758
rect -3351 -1078 3095 -842
rect 3331 -1078 3351 -842
rect -3351 -1162 3351 -1078
rect -3351 -1398 3095 -1162
rect 3331 -1398 3351 -1162
rect -3351 -1482 3351 -1398
rect -3351 -1718 3095 -1482
rect 3331 -1718 3351 -1482
rect -3351 -1802 3351 -1718
rect -3351 -2038 3095 -1802
rect 3331 -2038 3351 -1802
rect -3351 -2122 3351 -2038
rect -3351 -2358 3095 -2122
rect 3331 -2358 3351 -2122
rect -3351 -2442 3351 -2358
rect -3351 -2678 3095 -2442
rect 3331 -2678 3351 -2442
rect -3351 -2762 3351 -2678
rect -3351 -2998 3095 -2762
rect 3331 -2998 3351 -2762
rect -3351 -3100 3351 -2998
<< via4 >>
rect 3095 2762 3331 2998
rect 3095 2442 3331 2678
rect 3095 2122 3331 2358
rect 3095 1802 3331 2038
rect 3095 1482 3331 1718
rect 3095 1162 3331 1398
rect 3095 842 3331 1078
rect 3095 522 3331 758
rect 3095 202 3331 438
rect 3095 -118 3331 118
rect 3095 -438 3331 -202
rect 3095 -758 3331 -522
rect 3095 -1078 3331 -842
rect 3095 -1398 3331 -1162
rect 3095 -1718 3331 -1482
rect 3095 -2038 3331 -1802
rect 3095 -2358 3331 -2122
rect 3095 -2678 3331 -2442
rect 3095 -2998 3331 -2762
<< mimcap2 >>
rect -3251 2838 2749 3000
rect -3251 -2838 -3089 2838
rect 2587 -2838 2749 2838
rect -3251 -3000 2749 -2838
<< mimcap2contact >>
rect -3089 -2838 2587 2838
<< metal5 >>
rect 3053 2998 3373 3101
rect -3235 2838 2733 2984
rect -3235 -2838 -3089 2838
rect 2587 -2838 2733 2838
rect -3235 -2984 2733 -2838
rect 3053 2762 3095 2998
rect 3331 2762 3373 2998
rect 3053 2678 3373 2762
rect 3053 2442 3095 2678
rect 3331 2442 3373 2678
rect 3053 2358 3373 2442
rect 3053 2122 3095 2358
rect 3331 2122 3373 2358
rect 3053 2038 3373 2122
rect 3053 1802 3095 2038
rect 3331 1802 3373 2038
rect 3053 1718 3373 1802
rect 3053 1482 3095 1718
rect 3331 1482 3373 1718
rect 3053 1398 3373 1482
rect 3053 1162 3095 1398
rect 3331 1162 3373 1398
rect 3053 1078 3373 1162
rect 3053 842 3095 1078
rect 3331 842 3373 1078
rect 3053 758 3373 842
rect 3053 522 3095 758
rect 3331 522 3373 758
rect 3053 438 3373 522
rect 3053 202 3095 438
rect 3331 202 3373 438
rect 3053 118 3373 202
rect 3053 -118 3095 118
rect 3331 -118 3373 118
rect 3053 -202 3373 -118
rect 3053 -438 3095 -202
rect 3331 -438 3373 -202
rect 3053 -522 3373 -438
rect 3053 -758 3095 -522
rect 3331 -758 3373 -522
rect 3053 -842 3373 -758
rect 3053 -1078 3095 -842
rect 3331 -1078 3373 -842
rect 3053 -1162 3373 -1078
rect 3053 -1398 3095 -1162
rect 3331 -1398 3373 -1162
rect 3053 -1482 3373 -1398
rect 3053 -1718 3095 -1482
rect 3331 -1718 3373 -1482
rect 3053 -1802 3373 -1718
rect 3053 -2038 3095 -1802
rect 3331 -2038 3373 -1802
rect 3053 -2122 3373 -2038
rect 3053 -2358 3095 -2122
rect 3331 -2358 3373 -2122
rect 3053 -2442 3373 -2358
rect 3053 -2678 3095 -2442
rect 3331 -2678 3373 -2442
rect 3053 -2762 3373 -2678
rect 3053 -2998 3095 -2762
rect 3331 -2998 3373 -2762
rect 3053 -3101 3373 -2998
<< properties >>
string FIXED_BBOX -3351 -3100 2849 3100
<< end >>
