magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< error_p >>
rect -29 472 29 478
rect -29 438 -17 472
rect -29 432 29 438
rect -125 -438 -67 -432
rect 67 -438 125 -432
rect -125 -472 -113 -438
rect 67 -472 79 -438
rect -125 -478 -67 -472
rect 67 -478 125 -472
<< pwell >>
rect -301 -600 301 600
<< nmoslvt >>
rect -111 -400 -81 400
rect -15 -400 15 400
rect 81 -400 111 400
<< ndiff >>
rect -173 357 -111 400
rect -173 323 -161 357
rect -127 323 -111 357
rect -173 289 -111 323
rect -173 255 -161 289
rect -127 255 -111 289
rect -173 221 -111 255
rect -173 187 -161 221
rect -127 187 -111 221
rect -173 153 -111 187
rect -173 119 -161 153
rect -127 119 -111 153
rect -173 85 -111 119
rect -173 51 -161 85
rect -127 51 -111 85
rect -173 17 -111 51
rect -173 -17 -161 17
rect -127 -17 -111 17
rect -173 -51 -111 -17
rect -173 -85 -161 -51
rect -127 -85 -111 -51
rect -173 -119 -111 -85
rect -173 -153 -161 -119
rect -127 -153 -111 -119
rect -173 -187 -111 -153
rect -173 -221 -161 -187
rect -127 -221 -111 -187
rect -173 -255 -111 -221
rect -173 -289 -161 -255
rect -127 -289 -111 -255
rect -173 -323 -111 -289
rect -173 -357 -161 -323
rect -127 -357 -111 -323
rect -173 -400 -111 -357
rect -81 357 -15 400
rect -81 323 -65 357
rect -31 323 -15 357
rect -81 289 -15 323
rect -81 255 -65 289
rect -31 255 -15 289
rect -81 221 -15 255
rect -81 187 -65 221
rect -31 187 -15 221
rect -81 153 -15 187
rect -81 119 -65 153
rect -31 119 -15 153
rect -81 85 -15 119
rect -81 51 -65 85
rect -31 51 -15 85
rect -81 17 -15 51
rect -81 -17 -65 17
rect -31 -17 -15 17
rect -81 -51 -15 -17
rect -81 -85 -65 -51
rect -31 -85 -15 -51
rect -81 -119 -15 -85
rect -81 -153 -65 -119
rect -31 -153 -15 -119
rect -81 -187 -15 -153
rect -81 -221 -65 -187
rect -31 -221 -15 -187
rect -81 -255 -15 -221
rect -81 -289 -65 -255
rect -31 -289 -15 -255
rect -81 -323 -15 -289
rect -81 -357 -65 -323
rect -31 -357 -15 -323
rect -81 -400 -15 -357
rect 15 357 81 400
rect 15 323 31 357
rect 65 323 81 357
rect 15 289 81 323
rect 15 255 31 289
rect 65 255 81 289
rect 15 221 81 255
rect 15 187 31 221
rect 65 187 81 221
rect 15 153 81 187
rect 15 119 31 153
rect 65 119 81 153
rect 15 85 81 119
rect 15 51 31 85
rect 65 51 81 85
rect 15 17 81 51
rect 15 -17 31 17
rect 65 -17 81 17
rect 15 -51 81 -17
rect 15 -85 31 -51
rect 65 -85 81 -51
rect 15 -119 81 -85
rect 15 -153 31 -119
rect 65 -153 81 -119
rect 15 -187 81 -153
rect 15 -221 31 -187
rect 65 -221 81 -187
rect 15 -255 81 -221
rect 15 -289 31 -255
rect 65 -289 81 -255
rect 15 -323 81 -289
rect 15 -357 31 -323
rect 65 -357 81 -323
rect 15 -400 81 -357
rect 111 357 173 400
rect 111 323 127 357
rect 161 323 173 357
rect 111 289 173 323
rect 111 255 127 289
rect 161 255 173 289
rect 111 221 173 255
rect 111 187 127 221
rect 161 187 173 221
rect 111 153 173 187
rect 111 119 127 153
rect 161 119 173 153
rect 111 85 173 119
rect 111 51 127 85
rect 161 51 173 85
rect 111 17 173 51
rect 111 -17 127 17
rect 161 -17 173 17
rect 111 -51 173 -17
rect 111 -85 127 -51
rect 161 -85 173 -51
rect 111 -119 173 -85
rect 111 -153 127 -119
rect 161 -153 173 -119
rect 111 -187 173 -153
rect 111 -221 127 -187
rect 161 -221 173 -187
rect 111 -255 173 -221
rect 111 -289 127 -255
rect 161 -289 173 -255
rect 111 -323 173 -289
rect 111 -357 127 -323
rect 161 -357 173 -323
rect 111 -400 173 -357
<< ndiffc >>
rect -161 323 -127 357
rect -161 255 -127 289
rect -161 187 -127 221
rect -161 119 -127 153
rect -161 51 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -51
rect -161 -153 -127 -119
rect -161 -221 -127 -187
rect -161 -289 -127 -255
rect -161 -357 -127 -323
rect -65 323 -31 357
rect -65 255 -31 289
rect -65 187 -31 221
rect -65 119 -31 153
rect -65 51 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -51
rect -65 -153 -31 -119
rect -65 -221 -31 -187
rect -65 -289 -31 -255
rect -65 -357 -31 -323
rect 31 323 65 357
rect 31 255 65 289
rect 31 187 65 221
rect 31 119 65 153
rect 31 51 65 85
rect 31 -17 65 17
rect 31 -85 65 -51
rect 31 -153 65 -119
rect 31 -221 65 -187
rect 31 -289 65 -255
rect 31 -357 65 -323
rect 127 323 161 357
rect 127 255 161 289
rect 127 187 161 221
rect 127 119 161 153
rect 127 51 161 85
rect 127 -17 161 17
rect 127 -85 161 -51
rect 127 -153 161 -119
rect 127 -221 161 -187
rect 127 -289 161 -255
rect 127 -357 161 -323
<< psubdiff >>
rect -275 540 -153 574
rect -119 540 -85 574
rect -51 540 -17 574
rect 17 540 51 574
rect 85 540 119 574
rect 153 540 275 574
rect -275 459 -241 540
rect -275 391 -241 425
rect 241 459 275 540
rect -275 323 -241 357
rect -275 255 -241 289
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect -275 -289 -241 -255
rect -275 -357 -241 -323
rect -275 -425 -241 -391
rect 241 391 275 425
rect 241 323 275 357
rect 241 255 275 289
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect 241 -289 275 -255
rect 241 -357 275 -323
rect -275 -540 -241 -459
rect 241 -425 275 -391
rect 241 -540 275 -459
rect -275 -574 -153 -540
rect -119 -574 -85 -540
rect -51 -574 -17 -540
rect 17 -574 51 -540
rect 85 -574 119 -540
rect 153 -574 275 -540
<< psubdiffcont >>
rect -153 540 -119 574
rect -85 540 -51 574
rect -17 540 17 574
rect 51 540 85 574
rect 119 540 153 574
rect -275 425 -241 459
rect 241 425 275 459
rect -275 357 -241 391
rect -275 289 -241 323
rect -275 221 -241 255
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect -275 -255 -241 -221
rect -275 -323 -241 -289
rect -275 -391 -241 -357
rect 241 357 275 391
rect 241 289 275 323
rect 241 221 275 255
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect 241 -255 275 -221
rect 241 -323 275 -289
rect 241 -391 275 -357
rect -275 -459 -241 -425
rect 241 -459 275 -425
rect -153 -574 -119 -540
rect -85 -574 -51 -540
rect -17 -574 17 -540
rect 51 -574 85 -540
rect 119 -574 153 -540
<< poly >>
rect -33 472 33 488
rect -33 438 -17 472
rect 17 438 33 472
rect -111 400 -81 426
rect -33 422 33 438
rect -15 400 15 422
rect 81 400 111 426
rect -111 -422 -81 -400
rect -129 -438 -63 -422
rect -15 -426 15 -400
rect 81 -422 111 -400
rect -129 -472 -113 -438
rect -79 -472 -63 -438
rect -129 -488 -63 -472
rect 63 -438 129 -422
rect 63 -472 79 -438
rect 113 -472 129 -438
rect 63 -488 129 -472
<< polycont >>
rect -17 438 17 472
rect -113 -472 -79 -438
rect 79 -472 113 -438
<< locali >>
rect -275 540 -153 574
rect -119 540 -85 574
rect -51 540 -17 574
rect 17 540 51 574
rect 85 540 119 574
rect 153 540 275 574
rect -275 459 -241 540
rect -33 438 -17 472
rect 17 438 33 472
rect 241 459 275 540
rect -275 391 -241 425
rect -275 323 -241 357
rect -275 255 -241 289
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect -275 -289 -241 -255
rect -275 -357 -241 -323
rect -275 -425 -241 -391
rect -161 377 -127 404
rect -161 305 -127 323
rect -161 233 -127 255
rect -161 161 -127 187
rect -161 89 -127 119
rect -161 17 -127 51
rect -161 -51 -127 -17
rect -161 -119 -127 -89
rect -161 -187 -127 -161
rect -161 -255 -127 -233
rect -161 -323 -127 -305
rect -161 -404 -127 -377
rect -65 377 -31 404
rect -65 305 -31 323
rect -65 233 -31 255
rect -65 161 -31 187
rect -65 89 -31 119
rect -65 17 -31 51
rect -65 -51 -31 -17
rect -65 -119 -31 -89
rect -65 -187 -31 -161
rect -65 -255 -31 -233
rect -65 -323 -31 -305
rect -65 -404 -31 -377
rect 31 377 65 404
rect 31 305 65 323
rect 31 233 65 255
rect 31 161 65 187
rect 31 89 65 119
rect 31 17 65 51
rect 31 -51 65 -17
rect 31 -119 65 -89
rect 31 -187 65 -161
rect 31 -255 65 -233
rect 31 -323 65 -305
rect 31 -404 65 -377
rect 127 377 161 404
rect 127 305 161 323
rect 127 233 161 255
rect 127 161 161 187
rect 127 89 161 119
rect 127 17 161 51
rect 127 -51 161 -17
rect 127 -119 161 -89
rect 127 -187 161 -161
rect 127 -255 161 -233
rect 127 -323 161 -305
rect 127 -404 161 -377
rect 241 391 275 425
rect 241 323 275 357
rect 241 255 275 289
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect 241 -289 275 -255
rect 241 -357 275 -323
rect 241 -425 275 -391
rect -275 -540 -241 -459
rect -129 -472 -113 -438
rect -79 -472 -63 -438
rect 63 -472 79 -438
rect 113 -472 129 -438
rect 241 -540 275 -459
rect -275 -574 -153 -540
rect -119 -574 -85 -540
rect -51 -574 -17 -540
rect 17 -574 51 -540
rect 85 -574 119 -540
rect 153 -574 275 -540
<< viali >>
rect -17 438 17 472
rect -161 357 -127 377
rect -161 343 -127 357
rect -161 289 -127 305
rect -161 271 -127 289
rect -161 221 -127 233
rect -161 199 -127 221
rect -161 153 -127 161
rect -161 127 -127 153
rect -161 85 -127 89
rect -161 55 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -55
rect -161 -89 -127 -85
rect -161 -153 -127 -127
rect -161 -161 -127 -153
rect -161 -221 -127 -199
rect -161 -233 -127 -221
rect -161 -289 -127 -271
rect -161 -305 -127 -289
rect -161 -357 -127 -343
rect -161 -377 -127 -357
rect -65 357 -31 377
rect -65 343 -31 357
rect -65 289 -31 305
rect -65 271 -31 289
rect -65 221 -31 233
rect -65 199 -31 221
rect -65 153 -31 161
rect -65 127 -31 153
rect -65 85 -31 89
rect -65 55 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -55
rect -65 -89 -31 -85
rect -65 -153 -31 -127
rect -65 -161 -31 -153
rect -65 -221 -31 -199
rect -65 -233 -31 -221
rect -65 -289 -31 -271
rect -65 -305 -31 -289
rect -65 -357 -31 -343
rect -65 -377 -31 -357
rect 31 357 65 377
rect 31 343 65 357
rect 31 289 65 305
rect 31 271 65 289
rect 31 221 65 233
rect 31 199 65 221
rect 31 153 65 161
rect 31 127 65 153
rect 31 85 65 89
rect 31 55 65 85
rect 31 -17 65 17
rect 31 -85 65 -55
rect 31 -89 65 -85
rect 31 -153 65 -127
rect 31 -161 65 -153
rect 31 -221 65 -199
rect 31 -233 65 -221
rect 31 -289 65 -271
rect 31 -305 65 -289
rect 31 -357 65 -343
rect 31 -377 65 -357
rect 127 357 161 377
rect 127 343 161 357
rect 127 289 161 305
rect 127 271 161 289
rect 127 221 161 233
rect 127 199 161 221
rect 127 153 161 161
rect 127 127 161 153
rect 127 85 161 89
rect 127 55 161 85
rect 127 -17 161 17
rect 127 -85 161 -55
rect 127 -89 161 -85
rect 127 -153 161 -127
rect 127 -161 161 -153
rect 127 -221 161 -199
rect 127 -233 161 -221
rect 127 -289 161 -271
rect 127 -305 161 -289
rect 127 -357 161 -343
rect 127 -377 161 -357
rect -113 -472 -79 -438
rect 79 -472 113 -438
<< metal1 >>
rect -29 472 29 478
rect -29 438 -17 472
rect 17 438 29 472
rect -29 432 29 438
rect -167 377 -121 400
rect -167 343 -161 377
rect -127 343 -121 377
rect -167 305 -121 343
rect -167 271 -161 305
rect -127 271 -121 305
rect -167 233 -121 271
rect -167 199 -161 233
rect -127 199 -121 233
rect -167 161 -121 199
rect -167 127 -161 161
rect -127 127 -121 161
rect -167 89 -121 127
rect -167 55 -161 89
rect -127 55 -121 89
rect -167 17 -121 55
rect -167 -17 -161 17
rect -127 -17 -121 17
rect -167 -55 -121 -17
rect -167 -89 -161 -55
rect -127 -89 -121 -55
rect -167 -127 -121 -89
rect -167 -161 -161 -127
rect -127 -161 -121 -127
rect -167 -199 -121 -161
rect -167 -233 -161 -199
rect -127 -233 -121 -199
rect -167 -271 -121 -233
rect -167 -305 -161 -271
rect -127 -305 -121 -271
rect -167 -343 -121 -305
rect -167 -377 -161 -343
rect -127 -377 -121 -343
rect -167 -400 -121 -377
rect -71 377 -25 400
rect -71 343 -65 377
rect -31 343 -25 377
rect -71 305 -25 343
rect -71 271 -65 305
rect -31 271 -25 305
rect -71 233 -25 271
rect -71 199 -65 233
rect -31 199 -25 233
rect -71 161 -25 199
rect -71 127 -65 161
rect -31 127 -25 161
rect -71 89 -25 127
rect -71 55 -65 89
rect -31 55 -25 89
rect -71 17 -25 55
rect -71 -17 -65 17
rect -31 -17 -25 17
rect -71 -55 -25 -17
rect -71 -89 -65 -55
rect -31 -89 -25 -55
rect -71 -127 -25 -89
rect -71 -161 -65 -127
rect -31 -161 -25 -127
rect -71 -199 -25 -161
rect -71 -233 -65 -199
rect -31 -233 -25 -199
rect -71 -271 -25 -233
rect -71 -305 -65 -271
rect -31 -305 -25 -271
rect -71 -343 -25 -305
rect -71 -377 -65 -343
rect -31 -377 -25 -343
rect -71 -400 -25 -377
rect 25 377 71 400
rect 25 343 31 377
rect 65 343 71 377
rect 25 305 71 343
rect 25 271 31 305
rect 65 271 71 305
rect 25 233 71 271
rect 25 199 31 233
rect 65 199 71 233
rect 25 161 71 199
rect 25 127 31 161
rect 65 127 71 161
rect 25 89 71 127
rect 25 55 31 89
rect 65 55 71 89
rect 25 17 71 55
rect 25 -17 31 17
rect 65 -17 71 17
rect 25 -55 71 -17
rect 25 -89 31 -55
rect 65 -89 71 -55
rect 25 -127 71 -89
rect 25 -161 31 -127
rect 65 -161 71 -127
rect 25 -199 71 -161
rect 25 -233 31 -199
rect 65 -233 71 -199
rect 25 -271 71 -233
rect 25 -305 31 -271
rect 65 -305 71 -271
rect 25 -343 71 -305
rect 25 -377 31 -343
rect 65 -377 71 -343
rect 25 -400 71 -377
rect 121 377 167 400
rect 121 343 127 377
rect 161 343 167 377
rect 121 305 167 343
rect 121 271 127 305
rect 161 271 167 305
rect 121 233 167 271
rect 121 199 127 233
rect 161 199 167 233
rect 121 161 167 199
rect 121 127 127 161
rect 161 127 167 161
rect 121 89 167 127
rect 121 55 127 89
rect 161 55 167 89
rect 121 17 167 55
rect 121 -17 127 17
rect 161 -17 167 17
rect 121 -55 167 -17
rect 121 -89 127 -55
rect 161 -89 167 -55
rect 121 -127 167 -89
rect 121 -161 127 -127
rect 161 -161 167 -127
rect 121 -199 167 -161
rect 121 -233 127 -199
rect 161 -233 167 -199
rect 121 -271 167 -233
rect 121 -305 127 -271
rect 161 -305 167 -271
rect 121 -343 167 -305
rect 121 -377 127 -343
rect 161 -377 167 -343
rect 121 -400 167 -377
rect -125 -438 -67 -432
rect -125 -472 -113 -438
rect -79 -472 -67 -438
rect -125 -478 -67 -472
rect 67 -438 125 -432
rect 67 -472 79 -438
rect 113 -472 125 -438
rect 67 -478 125 -472
<< properties >>
string FIXED_BBOX -258 -557 258 557
<< end >>
