magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< metal4 >>
rect -2351 2038 2351 2100
rect -2351 1802 2095 2038
rect 2331 1802 2351 2038
rect -2351 1718 2351 1802
rect -2351 1482 2095 1718
rect 2331 1482 2351 1718
rect -2351 1398 2351 1482
rect -2351 1162 2095 1398
rect 2331 1162 2351 1398
rect -2351 1078 2351 1162
rect -2351 842 2095 1078
rect 2331 842 2351 1078
rect -2351 758 2351 842
rect -2351 522 2095 758
rect 2331 522 2351 758
rect -2351 438 2351 522
rect -2351 202 2095 438
rect 2331 202 2351 438
rect -2351 118 2351 202
rect -2351 -118 2095 118
rect 2331 -118 2351 118
rect -2351 -202 2351 -118
rect -2351 -438 2095 -202
rect 2331 -438 2351 -202
rect -2351 -522 2351 -438
rect -2351 -758 2095 -522
rect 2331 -758 2351 -522
rect -2351 -842 2351 -758
rect -2351 -1078 2095 -842
rect 2331 -1078 2351 -842
rect -2351 -1162 2351 -1078
rect -2351 -1398 2095 -1162
rect 2331 -1398 2351 -1162
rect -2351 -1482 2351 -1398
rect -2351 -1718 2095 -1482
rect 2331 -1718 2351 -1482
rect -2351 -1802 2351 -1718
rect -2351 -2038 2095 -1802
rect 2331 -2038 2351 -1802
rect -2351 -2100 2351 -2038
<< via4 >>
rect 2095 1802 2331 2038
rect 2095 1482 2331 1718
rect 2095 1162 2331 1398
rect 2095 842 2331 1078
rect 2095 522 2331 758
rect 2095 202 2331 438
rect 2095 -118 2331 118
rect 2095 -438 2331 -202
rect 2095 -758 2331 -522
rect 2095 -1078 2331 -842
rect 2095 -1398 2331 -1162
rect 2095 -1718 2331 -1482
rect 2095 -2038 2331 -1802
<< mimcap2 >>
rect -2251 1878 1749 2000
rect -2251 -1878 -2129 1878
rect 1627 -1878 1749 1878
rect -2251 -2000 1749 -1878
<< mimcap2contact >>
rect -2129 -1878 1627 1878
<< metal5 >>
rect 2053 2038 2373 2101
rect -2235 1878 1733 1984
rect -2235 -1878 -2129 1878
rect 1627 -1878 1733 1878
rect -2235 -1984 1733 -1878
rect 2053 1802 2095 2038
rect 2331 1802 2373 2038
rect 2053 1718 2373 1802
rect 2053 1482 2095 1718
rect 2331 1482 2373 1718
rect 2053 1398 2373 1482
rect 2053 1162 2095 1398
rect 2331 1162 2373 1398
rect 2053 1078 2373 1162
rect 2053 842 2095 1078
rect 2331 842 2373 1078
rect 2053 758 2373 842
rect 2053 522 2095 758
rect 2331 522 2373 758
rect 2053 438 2373 522
rect 2053 202 2095 438
rect 2331 202 2373 438
rect 2053 118 2373 202
rect 2053 -118 2095 118
rect 2331 -118 2373 118
rect 2053 -202 2373 -118
rect 2053 -438 2095 -202
rect 2331 -438 2373 -202
rect 2053 -522 2373 -438
rect 2053 -758 2095 -522
rect 2331 -758 2373 -522
rect 2053 -842 2373 -758
rect 2053 -1078 2095 -842
rect 2331 -1078 2373 -842
rect 2053 -1162 2373 -1078
rect 2053 -1398 2095 -1162
rect 2331 -1398 2373 -1162
rect 2053 -1482 2373 -1398
rect 2053 -1718 2095 -1482
rect 2331 -1718 2373 -1482
rect 2053 -1802 2373 -1718
rect 2053 -2038 2095 -1802
rect 2331 -2038 2373 -1802
rect 2053 -2101 2373 -2038
<< properties >>
string FIXED_BBOX -2351 -2100 1849 2100
<< end >>
