magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< error_p >>
rect -365 472 -307 478
rect -173 472 -115 478
rect 19 472 77 478
rect 211 472 269 478
rect 403 472 461 478
rect -365 438 -353 472
rect -173 438 -161 472
rect 19 438 31 472
rect 211 438 223 472
rect 403 438 415 472
rect -365 432 -307 438
rect -173 432 -115 438
rect 19 432 77 438
rect 211 432 269 438
rect 403 432 461 438
rect -461 -438 -403 -432
rect -269 -438 -211 -432
rect -77 -438 -19 -432
rect 115 -438 173 -432
rect 307 -438 365 -432
rect -461 -472 -449 -438
rect -269 -472 -257 -438
rect -77 -472 -65 -438
rect 115 -472 127 -438
rect 307 -472 319 -438
rect -461 -478 -403 -472
rect -269 -478 -211 -472
rect -77 -478 -19 -472
rect 115 -478 173 -472
rect 307 -478 365 -472
<< pwell >>
rect -637 -600 637 600
<< nmoslvt >>
rect -447 -400 -417 400
rect -351 -400 -321 400
rect -255 -400 -225 400
rect -159 -400 -129 400
rect -63 -400 -33 400
rect 33 -400 63 400
rect 129 -400 159 400
rect 225 -400 255 400
rect 321 -400 351 400
rect 417 -400 447 400
<< ndiff >>
rect -509 357 -447 400
rect -509 323 -497 357
rect -463 323 -447 357
rect -509 289 -447 323
rect -509 255 -497 289
rect -463 255 -447 289
rect -509 221 -447 255
rect -509 187 -497 221
rect -463 187 -447 221
rect -509 153 -447 187
rect -509 119 -497 153
rect -463 119 -447 153
rect -509 85 -447 119
rect -509 51 -497 85
rect -463 51 -447 85
rect -509 17 -447 51
rect -509 -17 -497 17
rect -463 -17 -447 17
rect -509 -51 -447 -17
rect -509 -85 -497 -51
rect -463 -85 -447 -51
rect -509 -119 -447 -85
rect -509 -153 -497 -119
rect -463 -153 -447 -119
rect -509 -187 -447 -153
rect -509 -221 -497 -187
rect -463 -221 -447 -187
rect -509 -255 -447 -221
rect -509 -289 -497 -255
rect -463 -289 -447 -255
rect -509 -323 -447 -289
rect -509 -357 -497 -323
rect -463 -357 -447 -323
rect -509 -400 -447 -357
rect -417 357 -351 400
rect -417 323 -401 357
rect -367 323 -351 357
rect -417 289 -351 323
rect -417 255 -401 289
rect -367 255 -351 289
rect -417 221 -351 255
rect -417 187 -401 221
rect -367 187 -351 221
rect -417 153 -351 187
rect -417 119 -401 153
rect -367 119 -351 153
rect -417 85 -351 119
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -119 -351 -85
rect -417 -153 -401 -119
rect -367 -153 -351 -119
rect -417 -187 -351 -153
rect -417 -221 -401 -187
rect -367 -221 -351 -187
rect -417 -255 -351 -221
rect -417 -289 -401 -255
rect -367 -289 -351 -255
rect -417 -323 -351 -289
rect -417 -357 -401 -323
rect -367 -357 -351 -323
rect -417 -400 -351 -357
rect -321 357 -255 400
rect -321 323 -305 357
rect -271 323 -255 357
rect -321 289 -255 323
rect -321 255 -305 289
rect -271 255 -255 289
rect -321 221 -255 255
rect -321 187 -305 221
rect -271 187 -255 221
rect -321 153 -255 187
rect -321 119 -305 153
rect -271 119 -255 153
rect -321 85 -255 119
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -119 -255 -85
rect -321 -153 -305 -119
rect -271 -153 -255 -119
rect -321 -187 -255 -153
rect -321 -221 -305 -187
rect -271 -221 -255 -187
rect -321 -255 -255 -221
rect -321 -289 -305 -255
rect -271 -289 -255 -255
rect -321 -323 -255 -289
rect -321 -357 -305 -323
rect -271 -357 -255 -323
rect -321 -400 -255 -357
rect -225 357 -159 400
rect -225 323 -209 357
rect -175 323 -159 357
rect -225 289 -159 323
rect -225 255 -209 289
rect -175 255 -159 289
rect -225 221 -159 255
rect -225 187 -209 221
rect -175 187 -159 221
rect -225 153 -159 187
rect -225 119 -209 153
rect -175 119 -159 153
rect -225 85 -159 119
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -119 -159 -85
rect -225 -153 -209 -119
rect -175 -153 -159 -119
rect -225 -187 -159 -153
rect -225 -221 -209 -187
rect -175 -221 -159 -187
rect -225 -255 -159 -221
rect -225 -289 -209 -255
rect -175 -289 -159 -255
rect -225 -323 -159 -289
rect -225 -357 -209 -323
rect -175 -357 -159 -323
rect -225 -400 -159 -357
rect -129 357 -63 400
rect -129 323 -113 357
rect -79 323 -63 357
rect -129 289 -63 323
rect -129 255 -113 289
rect -79 255 -63 289
rect -129 221 -63 255
rect -129 187 -113 221
rect -79 187 -63 221
rect -129 153 -63 187
rect -129 119 -113 153
rect -79 119 -63 153
rect -129 85 -63 119
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -119 -63 -85
rect -129 -153 -113 -119
rect -79 -153 -63 -119
rect -129 -187 -63 -153
rect -129 -221 -113 -187
rect -79 -221 -63 -187
rect -129 -255 -63 -221
rect -129 -289 -113 -255
rect -79 -289 -63 -255
rect -129 -323 -63 -289
rect -129 -357 -113 -323
rect -79 -357 -63 -323
rect -129 -400 -63 -357
rect -33 357 33 400
rect -33 323 -17 357
rect 17 323 33 357
rect -33 289 33 323
rect -33 255 -17 289
rect 17 255 33 289
rect -33 221 33 255
rect -33 187 -17 221
rect 17 187 33 221
rect -33 153 33 187
rect -33 119 -17 153
rect 17 119 33 153
rect -33 85 33 119
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -119 33 -85
rect -33 -153 -17 -119
rect 17 -153 33 -119
rect -33 -187 33 -153
rect -33 -221 -17 -187
rect 17 -221 33 -187
rect -33 -255 33 -221
rect -33 -289 -17 -255
rect 17 -289 33 -255
rect -33 -323 33 -289
rect -33 -357 -17 -323
rect 17 -357 33 -323
rect -33 -400 33 -357
rect 63 357 129 400
rect 63 323 79 357
rect 113 323 129 357
rect 63 289 129 323
rect 63 255 79 289
rect 113 255 129 289
rect 63 221 129 255
rect 63 187 79 221
rect 113 187 129 221
rect 63 153 129 187
rect 63 119 79 153
rect 113 119 129 153
rect 63 85 129 119
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -119 129 -85
rect 63 -153 79 -119
rect 113 -153 129 -119
rect 63 -187 129 -153
rect 63 -221 79 -187
rect 113 -221 129 -187
rect 63 -255 129 -221
rect 63 -289 79 -255
rect 113 -289 129 -255
rect 63 -323 129 -289
rect 63 -357 79 -323
rect 113 -357 129 -323
rect 63 -400 129 -357
rect 159 357 225 400
rect 159 323 175 357
rect 209 323 225 357
rect 159 289 225 323
rect 159 255 175 289
rect 209 255 225 289
rect 159 221 225 255
rect 159 187 175 221
rect 209 187 225 221
rect 159 153 225 187
rect 159 119 175 153
rect 209 119 225 153
rect 159 85 225 119
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -119 225 -85
rect 159 -153 175 -119
rect 209 -153 225 -119
rect 159 -187 225 -153
rect 159 -221 175 -187
rect 209 -221 225 -187
rect 159 -255 225 -221
rect 159 -289 175 -255
rect 209 -289 225 -255
rect 159 -323 225 -289
rect 159 -357 175 -323
rect 209 -357 225 -323
rect 159 -400 225 -357
rect 255 357 321 400
rect 255 323 271 357
rect 305 323 321 357
rect 255 289 321 323
rect 255 255 271 289
rect 305 255 321 289
rect 255 221 321 255
rect 255 187 271 221
rect 305 187 321 221
rect 255 153 321 187
rect 255 119 271 153
rect 305 119 321 153
rect 255 85 321 119
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -119 321 -85
rect 255 -153 271 -119
rect 305 -153 321 -119
rect 255 -187 321 -153
rect 255 -221 271 -187
rect 305 -221 321 -187
rect 255 -255 321 -221
rect 255 -289 271 -255
rect 305 -289 321 -255
rect 255 -323 321 -289
rect 255 -357 271 -323
rect 305 -357 321 -323
rect 255 -400 321 -357
rect 351 357 417 400
rect 351 323 367 357
rect 401 323 417 357
rect 351 289 417 323
rect 351 255 367 289
rect 401 255 417 289
rect 351 221 417 255
rect 351 187 367 221
rect 401 187 417 221
rect 351 153 417 187
rect 351 119 367 153
rect 401 119 417 153
rect 351 85 417 119
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -119 417 -85
rect 351 -153 367 -119
rect 401 -153 417 -119
rect 351 -187 417 -153
rect 351 -221 367 -187
rect 401 -221 417 -187
rect 351 -255 417 -221
rect 351 -289 367 -255
rect 401 -289 417 -255
rect 351 -323 417 -289
rect 351 -357 367 -323
rect 401 -357 417 -323
rect 351 -400 417 -357
rect 447 357 509 400
rect 447 323 463 357
rect 497 323 509 357
rect 447 289 509 323
rect 447 255 463 289
rect 497 255 509 289
rect 447 221 509 255
rect 447 187 463 221
rect 497 187 509 221
rect 447 153 509 187
rect 447 119 463 153
rect 497 119 509 153
rect 447 85 509 119
rect 447 51 463 85
rect 497 51 509 85
rect 447 17 509 51
rect 447 -17 463 17
rect 497 -17 509 17
rect 447 -51 509 -17
rect 447 -85 463 -51
rect 497 -85 509 -51
rect 447 -119 509 -85
rect 447 -153 463 -119
rect 497 -153 509 -119
rect 447 -187 509 -153
rect 447 -221 463 -187
rect 497 -221 509 -187
rect 447 -255 509 -221
rect 447 -289 463 -255
rect 497 -289 509 -255
rect 447 -323 509 -289
rect 447 -357 463 -323
rect 497 -357 509 -323
rect 447 -400 509 -357
<< ndiffc >>
rect -497 323 -463 357
rect -497 255 -463 289
rect -497 187 -463 221
rect -497 119 -463 153
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -497 -153 -463 -119
rect -497 -221 -463 -187
rect -497 -289 -463 -255
rect -497 -357 -463 -323
rect -401 323 -367 357
rect -401 255 -367 289
rect -401 187 -367 221
rect -401 119 -367 153
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -401 -153 -367 -119
rect -401 -221 -367 -187
rect -401 -289 -367 -255
rect -401 -357 -367 -323
rect -305 323 -271 357
rect -305 255 -271 289
rect -305 187 -271 221
rect -305 119 -271 153
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -305 -153 -271 -119
rect -305 -221 -271 -187
rect -305 -289 -271 -255
rect -305 -357 -271 -323
rect -209 323 -175 357
rect -209 255 -175 289
rect -209 187 -175 221
rect -209 119 -175 153
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -209 -153 -175 -119
rect -209 -221 -175 -187
rect -209 -289 -175 -255
rect -209 -357 -175 -323
rect -113 323 -79 357
rect -113 255 -79 289
rect -113 187 -79 221
rect -113 119 -79 153
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -113 -153 -79 -119
rect -113 -221 -79 -187
rect -113 -289 -79 -255
rect -113 -357 -79 -323
rect -17 323 17 357
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect -17 -357 17 -323
rect 79 323 113 357
rect 79 255 113 289
rect 79 187 113 221
rect 79 119 113 153
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 79 -153 113 -119
rect 79 -221 113 -187
rect 79 -289 113 -255
rect 79 -357 113 -323
rect 175 323 209 357
rect 175 255 209 289
rect 175 187 209 221
rect 175 119 209 153
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 175 -153 209 -119
rect 175 -221 209 -187
rect 175 -289 209 -255
rect 175 -357 209 -323
rect 271 323 305 357
rect 271 255 305 289
rect 271 187 305 221
rect 271 119 305 153
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 271 -153 305 -119
rect 271 -221 305 -187
rect 271 -289 305 -255
rect 271 -357 305 -323
rect 367 323 401 357
rect 367 255 401 289
rect 367 187 401 221
rect 367 119 401 153
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 367 -153 401 -119
rect 367 -221 401 -187
rect 367 -289 401 -255
rect 367 -357 401 -323
rect 463 323 497 357
rect 463 255 497 289
rect 463 187 497 221
rect 463 119 497 153
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 463 -153 497 -119
rect 463 -221 497 -187
rect 463 -289 497 -255
rect 463 -357 497 -323
<< psubdiff >>
rect -611 540 -493 574
rect -459 540 -425 574
rect -391 540 -357 574
rect -323 540 -289 574
rect -255 540 -221 574
rect -187 540 -153 574
rect -119 540 -85 574
rect -51 540 -17 574
rect 17 540 51 574
rect 85 540 119 574
rect 153 540 187 574
rect 221 540 255 574
rect 289 540 323 574
rect 357 540 391 574
rect 425 540 459 574
rect 493 540 611 574
rect -611 459 -577 540
rect -611 391 -577 425
rect 577 459 611 540
rect -611 323 -577 357
rect -611 255 -577 289
rect -611 187 -577 221
rect -611 119 -577 153
rect -611 51 -577 85
rect -611 -17 -577 17
rect -611 -85 -577 -51
rect -611 -153 -577 -119
rect -611 -221 -577 -187
rect -611 -289 -577 -255
rect -611 -357 -577 -323
rect -611 -425 -577 -391
rect 577 391 611 425
rect 577 323 611 357
rect 577 255 611 289
rect 577 187 611 221
rect 577 119 611 153
rect 577 51 611 85
rect 577 -17 611 17
rect 577 -85 611 -51
rect 577 -153 611 -119
rect 577 -221 611 -187
rect 577 -289 611 -255
rect 577 -357 611 -323
rect -611 -540 -577 -459
rect 577 -425 611 -391
rect 577 -540 611 -459
rect -611 -574 -493 -540
rect -459 -574 -425 -540
rect -391 -574 -357 -540
rect -323 -574 -289 -540
rect -255 -574 -221 -540
rect -187 -574 -153 -540
rect -119 -574 -85 -540
rect -51 -574 -17 -540
rect 17 -574 51 -540
rect 85 -574 119 -540
rect 153 -574 187 -540
rect 221 -574 255 -540
rect 289 -574 323 -540
rect 357 -574 391 -540
rect 425 -574 459 -540
rect 493 -574 611 -540
<< psubdiffcont >>
rect -493 540 -459 574
rect -425 540 -391 574
rect -357 540 -323 574
rect -289 540 -255 574
rect -221 540 -187 574
rect -153 540 -119 574
rect -85 540 -51 574
rect -17 540 17 574
rect 51 540 85 574
rect 119 540 153 574
rect 187 540 221 574
rect 255 540 289 574
rect 323 540 357 574
rect 391 540 425 574
rect 459 540 493 574
rect -611 425 -577 459
rect 577 425 611 459
rect -611 357 -577 391
rect -611 289 -577 323
rect -611 221 -577 255
rect -611 153 -577 187
rect -611 85 -577 119
rect -611 17 -577 51
rect -611 -51 -577 -17
rect -611 -119 -577 -85
rect -611 -187 -577 -153
rect -611 -255 -577 -221
rect -611 -323 -577 -289
rect -611 -391 -577 -357
rect 577 357 611 391
rect 577 289 611 323
rect 577 221 611 255
rect 577 153 611 187
rect 577 85 611 119
rect 577 17 611 51
rect 577 -51 611 -17
rect 577 -119 611 -85
rect 577 -187 611 -153
rect 577 -255 611 -221
rect 577 -323 611 -289
rect 577 -391 611 -357
rect -611 -459 -577 -425
rect 577 -459 611 -425
rect -493 -574 -459 -540
rect -425 -574 -391 -540
rect -357 -574 -323 -540
rect -289 -574 -255 -540
rect -221 -574 -187 -540
rect -153 -574 -119 -540
rect -85 -574 -51 -540
rect -17 -574 17 -540
rect 51 -574 85 -540
rect 119 -574 153 -540
rect 187 -574 221 -540
rect 255 -574 289 -540
rect 323 -574 357 -540
rect 391 -574 425 -540
rect 459 -574 493 -540
<< poly >>
rect -369 472 -303 488
rect -369 438 -353 472
rect -319 438 -303 472
rect -447 400 -417 426
rect -369 422 -303 438
rect -177 472 -111 488
rect -177 438 -161 472
rect -127 438 -111 472
rect -351 400 -321 422
rect -255 400 -225 426
rect -177 422 -111 438
rect 15 472 81 488
rect 15 438 31 472
rect 65 438 81 472
rect -159 400 -129 422
rect -63 400 -33 426
rect 15 422 81 438
rect 207 472 273 488
rect 207 438 223 472
rect 257 438 273 472
rect 33 400 63 422
rect 129 400 159 426
rect 207 422 273 438
rect 399 472 465 488
rect 399 438 415 472
rect 449 438 465 472
rect 225 400 255 422
rect 321 400 351 426
rect 399 422 465 438
rect 417 400 447 422
rect -447 -422 -417 -400
rect -465 -438 -399 -422
rect -351 -426 -321 -400
rect -255 -422 -225 -400
rect -465 -472 -449 -438
rect -415 -472 -399 -438
rect -465 -488 -399 -472
rect -273 -438 -207 -422
rect -159 -426 -129 -400
rect -63 -422 -33 -400
rect -273 -472 -257 -438
rect -223 -472 -207 -438
rect -273 -488 -207 -472
rect -81 -438 -15 -422
rect 33 -426 63 -400
rect 129 -422 159 -400
rect -81 -472 -65 -438
rect -31 -472 -15 -438
rect -81 -488 -15 -472
rect 111 -438 177 -422
rect 225 -426 255 -400
rect 321 -422 351 -400
rect 111 -472 127 -438
rect 161 -472 177 -438
rect 111 -488 177 -472
rect 303 -438 369 -422
rect 417 -426 447 -400
rect 303 -472 319 -438
rect 353 -472 369 -438
rect 303 -488 369 -472
<< polycont >>
rect -353 438 -319 472
rect -161 438 -127 472
rect 31 438 65 472
rect 223 438 257 472
rect 415 438 449 472
rect -449 -472 -415 -438
rect -257 -472 -223 -438
rect -65 -472 -31 -438
rect 127 -472 161 -438
rect 319 -472 353 -438
<< locali >>
rect -611 540 -493 574
rect -459 540 -425 574
rect -391 540 -357 574
rect -323 540 -289 574
rect -255 540 -221 574
rect -187 540 -153 574
rect -119 540 -85 574
rect -51 540 -17 574
rect 17 540 51 574
rect 85 540 119 574
rect 153 540 187 574
rect 221 540 255 574
rect 289 540 323 574
rect 357 540 391 574
rect 425 540 459 574
rect 493 540 611 574
rect -611 459 -577 540
rect -369 438 -353 472
rect -319 438 -303 472
rect -177 438 -161 472
rect -127 438 -111 472
rect 15 438 31 472
rect 65 438 81 472
rect 207 438 223 472
rect 257 438 273 472
rect 399 438 415 472
rect 449 438 465 472
rect 577 459 611 540
rect -611 391 -577 425
rect -611 323 -577 357
rect -611 255 -577 289
rect -611 187 -577 221
rect -611 119 -577 153
rect -611 51 -577 85
rect -611 -17 -577 17
rect -611 -85 -577 -51
rect -611 -153 -577 -119
rect -611 -221 -577 -187
rect -611 -289 -577 -255
rect -611 -357 -577 -323
rect -611 -425 -577 -391
rect -497 377 -463 404
rect -497 305 -463 323
rect -497 233 -463 255
rect -497 161 -463 187
rect -497 89 -463 119
rect -497 17 -463 51
rect -497 -51 -463 -17
rect -497 -119 -463 -89
rect -497 -187 -463 -161
rect -497 -255 -463 -233
rect -497 -323 -463 -305
rect -497 -404 -463 -377
rect -401 377 -367 404
rect -401 305 -367 323
rect -401 233 -367 255
rect -401 161 -367 187
rect -401 89 -367 119
rect -401 17 -367 51
rect -401 -51 -367 -17
rect -401 -119 -367 -89
rect -401 -187 -367 -161
rect -401 -255 -367 -233
rect -401 -323 -367 -305
rect -401 -404 -367 -377
rect -305 377 -271 404
rect -305 305 -271 323
rect -305 233 -271 255
rect -305 161 -271 187
rect -305 89 -271 119
rect -305 17 -271 51
rect -305 -51 -271 -17
rect -305 -119 -271 -89
rect -305 -187 -271 -161
rect -305 -255 -271 -233
rect -305 -323 -271 -305
rect -305 -404 -271 -377
rect -209 377 -175 404
rect -209 305 -175 323
rect -209 233 -175 255
rect -209 161 -175 187
rect -209 89 -175 119
rect -209 17 -175 51
rect -209 -51 -175 -17
rect -209 -119 -175 -89
rect -209 -187 -175 -161
rect -209 -255 -175 -233
rect -209 -323 -175 -305
rect -209 -404 -175 -377
rect -113 377 -79 404
rect -113 305 -79 323
rect -113 233 -79 255
rect -113 161 -79 187
rect -113 89 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -89
rect -113 -187 -79 -161
rect -113 -255 -79 -233
rect -113 -323 -79 -305
rect -113 -404 -79 -377
rect -17 377 17 404
rect -17 305 17 323
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -323 17 -305
rect -17 -404 17 -377
rect 79 377 113 404
rect 79 305 113 323
rect 79 233 113 255
rect 79 161 113 187
rect 79 89 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -89
rect 79 -187 113 -161
rect 79 -255 113 -233
rect 79 -323 113 -305
rect 79 -404 113 -377
rect 175 377 209 404
rect 175 305 209 323
rect 175 233 209 255
rect 175 161 209 187
rect 175 89 209 119
rect 175 17 209 51
rect 175 -51 209 -17
rect 175 -119 209 -89
rect 175 -187 209 -161
rect 175 -255 209 -233
rect 175 -323 209 -305
rect 175 -404 209 -377
rect 271 377 305 404
rect 271 305 305 323
rect 271 233 305 255
rect 271 161 305 187
rect 271 89 305 119
rect 271 17 305 51
rect 271 -51 305 -17
rect 271 -119 305 -89
rect 271 -187 305 -161
rect 271 -255 305 -233
rect 271 -323 305 -305
rect 271 -404 305 -377
rect 367 377 401 404
rect 367 305 401 323
rect 367 233 401 255
rect 367 161 401 187
rect 367 89 401 119
rect 367 17 401 51
rect 367 -51 401 -17
rect 367 -119 401 -89
rect 367 -187 401 -161
rect 367 -255 401 -233
rect 367 -323 401 -305
rect 367 -404 401 -377
rect 463 377 497 404
rect 463 305 497 323
rect 463 233 497 255
rect 463 161 497 187
rect 463 89 497 119
rect 463 17 497 51
rect 463 -51 497 -17
rect 463 -119 497 -89
rect 463 -187 497 -161
rect 463 -255 497 -233
rect 463 -323 497 -305
rect 463 -404 497 -377
rect 577 391 611 425
rect 577 323 611 357
rect 577 255 611 289
rect 577 187 611 221
rect 577 119 611 153
rect 577 51 611 85
rect 577 -17 611 17
rect 577 -85 611 -51
rect 577 -153 611 -119
rect 577 -221 611 -187
rect 577 -289 611 -255
rect 577 -357 611 -323
rect 577 -425 611 -391
rect -611 -540 -577 -459
rect -465 -472 -449 -438
rect -415 -472 -399 -438
rect -273 -472 -257 -438
rect -223 -472 -207 -438
rect -81 -472 -65 -438
rect -31 -472 -15 -438
rect 111 -472 127 -438
rect 161 -472 177 -438
rect 303 -472 319 -438
rect 353 -472 369 -438
rect 577 -540 611 -459
rect -611 -574 -493 -540
rect -459 -574 -425 -540
rect -391 -574 -357 -540
rect -323 -574 -289 -540
rect -255 -574 -221 -540
rect -187 -574 -153 -540
rect -119 -574 -85 -540
rect -51 -574 -17 -540
rect 17 -574 51 -540
rect 85 -574 119 -540
rect 153 -574 187 -540
rect 221 -574 255 -540
rect 289 -574 323 -540
rect 357 -574 391 -540
rect 425 -574 459 -540
rect 493 -574 611 -540
<< viali >>
rect -353 438 -319 472
rect -161 438 -127 472
rect 31 438 65 472
rect 223 438 257 472
rect 415 438 449 472
rect -497 357 -463 377
rect -497 343 -463 357
rect -497 289 -463 305
rect -497 271 -463 289
rect -497 221 -463 233
rect -497 199 -463 221
rect -497 153 -463 161
rect -497 127 -463 153
rect -497 85 -463 89
rect -497 55 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -55
rect -497 -89 -463 -85
rect -497 -153 -463 -127
rect -497 -161 -463 -153
rect -497 -221 -463 -199
rect -497 -233 -463 -221
rect -497 -289 -463 -271
rect -497 -305 -463 -289
rect -497 -357 -463 -343
rect -497 -377 -463 -357
rect -401 357 -367 377
rect -401 343 -367 357
rect -401 289 -367 305
rect -401 271 -367 289
rect -401 221 -367 233
rect -401 199 -367 221
rect -401 153 -367 161
rect -401 127 -367 153
rect -401 85 -367 89
rect -401 55 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -55
rect -401 -89 -367 -85
rect -401 -153 -367 -127
rect -401 -161 -367 -153
rect -401 -221 -367 -199
rect -401 -233 -367 -221
rect -401 -289 -367 -271
rect -401 -305 -367 -289
rect -401 -357 -367 -343
rect -401 -377 -367 -357
rect -305 357 -271 377
rect -305 343 -271 357
rect -305 289 -271 305
rect -305 271 -271 289
rect -305 221 -271 233
rect -305 199 -271 221
rect -305 153 -271 161
rect -305 127 -271 153
rect -305 85 -271 89
rect -305 55 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -55
rect -305 -89 -271 -85
rect -305 -153 -271 -127
rect -305 -161 -271 -153
rect -305 -221 -271 -199
rect -305 -233 -271 -221
rect -305 -289 -271 -271
rect -305 -305 -271 -289
rect -305 -357 -271 -343
rect -305 -377 -271 -357
rect -209 357 -175 377
rect -209 343 -175 357
rect -209 289 -175 305
rect -209 271 -175 289
rect -209 221 -175 233
rect -209 199 -175 221
rect -209 153 -175 161
rect -209 127 -175 153
rect -209 85 -175 89
rect -209 55 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -55
rect -209 -89 -175 -85
rect -209 -153 -175 -127
rect -209 -161 -175 -153
rect -209 -221 -175 -199
rect -209 -233 -175 -221
rect -209 -289 -175 -271
rect -209 -305 -175 -289
rect -209 -357 -175 -343
rect -209 -377 -175 -357
rect -113 357 -79 377
rect -113 343 -79 357
rect -113 289 -79 305
rect -113 271 -79 289
rect -113 221 -79 233
rect -113 199 -79 221
rect -113 153 -79 161
rect -113 127 -79 153
rect -113 85 -79 89
rect -113 55 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -55
rect -113 -89 -79 -85
rect -113 -153 -79 -127
rect -113 -161 -79 -153
rect -113 -221 -79 -199
rect -113 -233 -79 -221
rect -113 -289 -79 -271
rect -113 -305 -79 -289
rect -113 -357 -79 -343
rect -113 -377 -79 -357
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect 79 357 113 377
rect 79 343 113 357
rect 79 289 113 305
rect 79 271 113 289
rect 79 221 113 233
rect 79 199 113 221
rect 79 153 113 161
rect 79 127 113 153
rect 79 85 113 89
rect 79 55 113 85
rect 79 -17 113 17
rect 79 -85 113 -55
rect 79 -89 113 -85
rect 79 -153 113 -127
rect 79 -161 113 -153
rect 79 -221 113 -199
rect 79 -233 113 -221
rect 79 -289 113 -271
rect 79 -305 113 -289
rect 79 -357 113 -343
rect 79 -377 113 -357
rect 175 357 209 377
rect 175 343 209 357
rect 175 289 209 305
rect 175 271 209 289
rect 175 221 209 233
rect 175 199 209 221
rect 175 153 209 161
rect 175 127 209 153
rect 175 85 209 89
rect 175 55 209 85
rect 175 -17 209 17
rect 175 -85 209 -55
rect 175 -89 209 -85
rect 175 -153 209 -127
rect 175 -161 209 -153
rect 175 -221 209 -199
rect 175 -233 209 -221
rect 175 -289 209 -271
rect 175 -305 209 -289
rect 175 -357 209 -343
rect 175 -377 209 -357
rect 271 357 305 377
rect 271 343 305 357
rect 271 289 305 305
rect 271 271 305 289
rect 271 221 305 233
rect 271 199 305 221
rect 271 153 305 161
rect 271 127 305 153
rect 271 85 305 89
rect 271 55 305 85
rect 271 -17 305 17
rect 271 -85 305 -55
rect 271 -89 305 -85
rect 271 -153 305 -127
rect 271 -161 305 -153
rect 271 -221 305 -199
rect 271 -233 305 -221
rect 271 -289 305 -271
rect 271 -305 305 -289
rect 271 -357 305 -343
rect 271 -377 305 -357
rect 367 357 401 377
rect 367 343 401 357
rect 367 289 401 305
rect 367 271 401 289
rect 367 221 401 233
rect 367 199 401 221
rect 367 153 401 161
rect 367 127 401 153
rect 367 85 401 89
rect 367 55 401 85
rect 367 -17 401 17
rect 367 -85 401 -55
rect 367 -89 401 -85
rect 367 -153 401 -127
rect 367 -161 401 -153
rect 367 -221 401 -199
rect 367 -233 401 -221
rect 367 -289 401 -271
rect 367 -305 401 -289
rect 367 -357 401 -343
rect 367 -377 401 -357
rect 463 357 497 377
rect 463 343 497 357
rect 463 289 497 305
rect 463 271 497 289
rect 463 221 497 233
rect 463 199 497 221
rect 463 153 497 161
rect 463 127 497 153
rect 463 85 497 89
rect 463 55 497 85
rect 463 -17 497 17
rect 463 -85 497 -55
rect 463 -89 497 -85
rect 463 -153 497 -127
rect 463 -161 497 -153
rect 463 -221 497 -199
rect 463 -233 497 -221
rect 463 -289 497 -271
rect 463 -305 497 -289
rect 463 -357 497 -343
rect 463 -377 497 -357
rect -449 -472 -415 -438
rect -257 -472 -223 -438
rect -65 -472 -31 -438
rect 127 -472 161 -438
rect 319 -472 353 -438
<< metal1 >>
rect -365 472 -307 478
rect -365 438 -353 472
rect -319 438 -307 472
rect -365 432 -307 438
rect -173 472 -115 478
rect -173 438 -161 472
rect -127 438 -115 472
rect -173 432 -115 438
rect 19 472 77 478
rect 19 438 31 472
rect 65 438 77 472
rect 19 432 77 438
rect 211 472 269 478
rect 211 438 223 472
rect 257 438 269 472
rect 211 432 269 438
rect 403 472 461 478
rect 403 438 415 472
rect 449 438 461 472
rect 403 432 461 438
rect -503 377 -457 400
rect -503 343 -497 377
rect -463 343 -457 377
rect -503 305 -457 343
rect -503 271 -497 305
rect -463 271 -457 305
rect -503 233 -457 271
rect -503 199 -497 233
rect -463 199 -457 233
rect -503 161 -457 199
rect -503 127 -497 161
rect -463 127 -457 161
rect -503 89 -457 127
rect -503 55 -497 89
rect -463 55 -457 89
rect -503 17 -457 55
rect -503 -17 -497 17
rect -463 -17 -457 17
rect -503 -55 -457 -17
rect -503 -89 -497 -55
rect -463 -89 -457 -55
rect -503 -127 -457 -89
rect -503 -161 -497 -127
rect -463 -161 -457 -127
rect -503 -199 -457 -161
rect -503 -233 -497 -199
rect -463 -233 -457 -199
rect -503 -271 -457 -233
rect -503 -305 -497 -271
rect -463 -305 -457 -271
rect -503 -343 -457 -305
rect -503 -377 -497 -343
rect -463 -377 -457 -343
rect -503 -400 -457 -377
rect -407 377 -361 400
rect -407 343 -401 377
rect -367 343 -361 377
rect -407 305 -361 343
rect -407 271 -401 305
rect -367 271 -361 305
rect -407 233 -361 271
rect -407 199 -401 233
rect -367 199 -361 233
rect -407 161 -361 199
rect -407 127 -401 161
rect -367 127 -361 161
rect -407 89 -361 127
rect -407 55 -401 89
rect -367 55 -361 89
rect -407 17 -361 55
rect -407 -17 -401 17
rect -367 -17 -361 17
rect -407 -55 -361 -17
rect -407 -89 -401 -55
rect -367 -89 -361 -55
rect -407 -127 -361 -89
rect -407 -161 -401 -127
rect -367 -161 -361 -127
rect -407 -199 -361 -161
rect -407 -233 -401 -199
rect -367 -233 -361 -199
rect -407 -271 -361 -233
rect -407 -305 -401 -271
rect -367 -305 -361 -271
rect -407 -343 -361 -305
rect -407 -377 -401 -343
rect -367 -377 -361 -343
rect -407 -400 -361 -377
rect -311 377 -265 400
rect -311 343 -305 377
rect -271 343 -265 377
rect -311 305 -265 343
rect -311 271 -305 305
rect -271 271 -265 305
rect -311 233 -265 271
rect -311 199 -305 233
rect -271 199 -265 233
rect -311 161 -265 199
rect -311 127 -305 161
rect -271 127 -265 161
rect -311 89 -265 127
rect -311 55 -305 89
rect -271 55 -265 89
rect -311 17 -265 55
rect -311 -17 -305 17
rect -271 -17 -265 17
rect -311 -55 -265 -17
rect -311 -89 -305 -55
rect -271 -89 -265 -55
rect -311 -127 -265 -89
rect -311 -161 -305 -127
rect -271 -161 -265 -127
rect -311 -199 -265 -161
rect -311 -233 -305 -199
rect -271 -233 -265 -199
rect -311 -271 -265 -233
rect -311 -305 -305 -271
rect -271 -305 -265 -271
rect -311 -343 -265 -305
rect -311 -377 -305 -343
rect -271 -377 -265 -343
rect -311 -400 -265 -377
rect -215 377 -169 400
rect -215 343 -209 377
rect -175 343 -169 377
rect -215 305 -169 343
rect -215 271 -209 305
rect -175 271 -169 305
rect -215 233 -169 271
rect -215 199 -209 233
rect -175 199 -169 233
rect -215 161 -169 199
rect -215 127 -209 161
rect -175 127 -169 161
rect -215 89 -169 127
rect -215 55 -209 89
rect -175 55 -169 89
rect -215 17 -169 55
rect -215 -17 -209 17
rect -175 -17 -169 17
rect -215 -55 -169 -17
rect -215 -89 -209 -55
rect -175 -89 -169 -55
rect -215 -127 -169 -89
rect -215 -161 -209 -127
rect -175 -161 -169 -127
rect -215 -199 -169 -161
rect -215 -233 -209 -199
rect -175 -233 -169 -199
rect -215 -271 -169 -233
rect -215 -305 -209 -271
rect -175 -305 -169 -271
rect -215 -343 -169 -305
rect -215 -377 -209 -343
rect -175 -377 -169 -343
rect -215 -400 -169 -377
rect -119 377 -73 400
rect -119 343 -113 377
rect -79 343 -73 377
rect -119 305 -73 343
rect -119 271 -113 305
rect -79 271 -73 305
rect -119 233 -73 271
rect -119 199 -113 233
rect -79 199 -73 233
rect -119 161 -73 199
rect -119 127 -113 161
rect -79 127 -73 161
rect -119 89 -73 127
rect -119 55 -113 89
rect -79 55 -73 89
rect -119 17 -73 55
rect -119 -17 -113 17
rect -79 -17 -73 17
rect -119 -55 -73 -17
rect -119 -89 -113 -55
rect -79 -89 -73 -55
rect -119 -127 -73 -89
rect -119 -161 -113 -127
rect -79 -161 -73 -127
rect -119 -199 -73 -161
rect -119 -233 -113 -199
rect -79 -233 -73 -199
rect -119 -271 -73 -233
rect -119 -305 -113 -271
rect -79 -305 -73 -271
rect -119 -343 -73 -305
rect -119 -377 -113 -343
rect -79 -377 -73 -343
rect -119 -400 -73 -377
rect -23 377 23 400
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -400 23 -377
rect 73 377 119 400
rect 73 343 79 377
rect 113 343 119 377
rect 73 305 119 343
rect 73 271 79 305
rect 113 271 119 305
rect 73 233 119 271
rect 73 199 79 233
rect 113 199 119 233
rect 73 161 119 199
rect 73 127 79 161
rect 113 127 119 161
rect 73 89 119 127
rect 73 55 79 89
rect 113 55 119 89
rect 73 17 119 55
rect 73 -17 79 17
rect 113 -17 119 17
rect 73 -55 119 -17
rect 73 -89 79 -55
rect 113 -89 119 -55
rect 73 -127 119 -89
rect 73 -161 79 -127
rect 113 -161 119 -127
rect 73 -199 119 -161
rect 73 -233 79 -199
rect 113 -233 119 -199
rect 73 -271 119 -233
rect 73 -305 79 -271
rect 113 -305 119 -271
rect 73 -343 119 -305
rect 73 -377 79 -343
rect 113 -377 119 -343
rect 73 -400 119 -377
rect 169 377 215 400
rect 169 343 175 377
rect 209 343 215 377
rect 169 305 215 343
rect 169 271 175 305
rect 209 271 215 305
rect 169 233 215 271
rect 169 199 175 233
rect 209 199 215 233
rect 169 161 215 199
rect 169 127 175 161
rect 209 127 215 161
rect 169 89 215 127
rect 169 55 175 89
rect 209 55 215 89
rect 169 17 215 55
rect 169 -17 175 17
rect 209 -17 215 17
rect 169 -55 215 -17
rect 169 -89 175 -55
rect 209 -89 215 -55
rect 169 -127 215 -89
rect 169 -161 175 -127
rect 209 -161 215 -127
rect 169 -199 215 -161
rect 169 -233 175 -199
rect 209 -233 215 -199
rect 169 -271 215 -233
rect 169 -305 175 -271
rect 209 -305 215 -271
rect 169 -343 215 -305
rect 169 -377 175 -343
rect 209 -377 215 -343
rect 169 -400 215 -377
rect 265 377 311 400
rect 265 343 271 377
rect 305 343 311 377
rect 265 305 311 343
rect 265 271 271 305
rect 305 271 311 305
rect 265 233 311 271
rect 265 199 271 233
rect 305 199 311 233
rect 265 161 311 199
rect 265 127 271 161
rect 305 127 311 161
rect 265 89 311 127
rect 265 55 271 89
rect 305 55 311 89
rect 265 17 311 55
rect 265 -17 271 17
rect 305 -17 311 17
rect 265 -55 311 -17
rect 265 -89 271 -55
rect 305 -89 311 -55
rect 265 -127 311 -89
rect 265 -161 271 -127
rect 305 -161 311 -127
rect 265 -199 311 -161
rect 265 -233 271 -199
rect 305 -233 311 -199
rect 265 -271 311 -233
rect 265 -305 271 -271
rect 305 -305 311 -271
rect 265 -343 311 -305
rect 265 -377 271 -343
rect 305 -377 311 -343
rect 265 -400 311 -377
rect 361 377 407 400
rect 361 343 367 377
rect 401 343 407 377
rect 361 305 407 343
rect 361 271 367 305
rect 401 271 407 305
rect 361 233 407 271
rect 361 199 367 233
rect 401 199 407 233
rect 361 161 407 199
rect 361 127 367 161
rect 401 127 407 161
rect 361 89 407 127
rect 361 55 367 89
rect 401 55 407 89
rect 361 17 407 55
rect 361 -17 367 17
rect 401 -17 407 17
rect 361 -55 407 -17
rect 361 -89 367 -55
rect 401 -89 407 -55
rect 361 -127 407 -89
rect 361 -161 367 -127
rect 401 -161 407 -127
rect 361 -199 407 -161
rect 361 -233 367 -199
rect 401 -233 407 -199
rect 361 -271 407 -233
rect 361 -305 367 -271
rect 401 -305 407 -271
rect 361 -343 407 -305
rect 361 -377 367 -343
rect 401 -377 407 -343
rect 361 -400 407 -377
rect 457 377 503 400
rect 457 343 463 377
rect 497 343 503 377
rect 457 305 503 343
rect 457 271 463 305
rect 497 271 503 305
rect 457 233 503 271
rect 457 199 463 233
rect 497 199 503 233
rect 457 161 503 199
rect 457 127 463 161
rect 497 127 503 161
rect 457 89 503 127
rect 457 55 463 89
rect 497 55 503 89
rect 457 17 503 55
rect 457 -17 463 17
rect 497 -17 503 17
rect 457 -55 503 -17
rect 457 -89 463 -55
rect 497 -89 503 -55
rect 457 -127 503 -89
rect 457 -161 463 -127
rect 497 -161 503 -127
rect 457 -199 503 -161
rect 457 -233 463 -199
rect 497 -233 503 -199
rect 457 -271 503 -233
rect 457 -305 463 -271
rect 497 -305 503 -271
rect 457 -343 503 -305
rect 457 -377 463 -343
rect 497 -377 503 -343
rect 457 -400 503 -377
rect -461 -438 -403 -432
rect -461 -472 -449 -438
rect -415 -472 -403 -438
rect -461 -478 -403 -472
rect -269 -438 -211 -432
rect -269 -472 -257 -438
rect -223 -472 -211 -438
rect -269 -478 -211 -472
rect -77 -438 -19 -432
rect -77 -472 -65 -438
rect -31 -472 -19 -438
rect -77 -478 -19 -472
rect 115 -438 173 -432
rect 115 -472 127 -438
rect 161 -472 173 -438
rect 115 -478 173 -472
rect 307 -438 365 -432
rect 307 -472 319 -438
rect 353 -472 365 -438
rect 307 -478 365 -472
<< properties >>
string FIXED_BBOX -594 -557 594 557
<< end >>
