magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< pwell >>
rect -804 571 804 657
rect -804 -571 -718 571
rect 718 -571 804 571
rect -804 -657 804 -571
<< psubdiff >>
rect -778 597 -663 631
rect -629 597 -595 631
rect -561 597 -527 631
rect -493 597 -459 631
rect -425 597 -391 631
rect -357 597 -323 631
rect -289 597 -255 631
rect -221 597 -187 631
rect -153 597 -119 631
rect -85 597 -51 631
rect -17 597 17 631
rect 51 597 85 631
rect 119 597 153 631
rect 187 597 221 631
rect 255 597 289 631
rect 323 597 357 631
rect 391 597 425 631
rect 459 597 493 631
rect 527 597 561 631
rect 595 597 629 631
rect 663 597 778 631
rect -778 527 -744 597
rect 744 527 778 597
rect -778 459 -744 493
rect -778 391 -744 425
rect -778 323 -744 357
rect -778 255 -744 289
rect -778 187 -744 221
rect -778 119 -744 153
rect -778 51 -744 85
rect -778 -17 -744 17
rect -778 -85 -744 -51
rect -778 -153 -744 -119
rect -778 -221 -744 -187
rect -778 -289 -744 -255
rect -778 -357 -744 -323
rect -778 -425 -744 -391
rect -778 -493 -744 -459
rect 744 459 778 493
rect 744 391 778 425
rect 744 323 778 357
rect 744 255 778 289
rect 744 187 778 221
rect 744 119 778 153
rect 744 51 778 85
rect 744 -17 778 17
rect 744 -85 778 -51
rect 744 -153 778 -119
rect 744 -221 778 -187
rect 744 -289 778 -255
rect 744 -357 778 -323
rect 744 -425 778 -391
rect 744 -493 778 -459
rect -778 -597 -744 -527
rect 744 -597 778 -527
rect -778 -631 -663 -597
rect -629 -631 -595 -597
rect -561 -631 -527 -597
rect -493 -631 -459 -597
rect -425 -631 -391 -597
rect -357 -631 -323 -597
rect -289 -631 -255 -597
rect -221 -631 -187 -597
rect -153 -631 -119 -597
rect -85 -631 -51 -597
rect -17 -631 17 -597
rect 51 -631 85 -597
rect 119 -631 153 -597
rect 187 -631 221 -597
rect 255 -631 289 -597
rect 323 -631 357 -597
rect 391 -631 425 -597
rect 459 -631 493 -597
rect 527 -631 561 -597
rect 595 -631 629 -597
rect 663 -631 778 -597
<< psubdiffcont >>
rect -663 597 -629 631
rect -595 597 -561 631
rect -527 597 -493 631
rect -459 597 -425 631
rect -391 597 -357 631
rect -323 597 -289 631
rect -255 597 -221 631
rect -187 597 -153 631
rect -119 597 -85 631
rect -51 597 -17 631
rect 17 597 51 631
rect 85 597 119 631
rect 153 597 187 631
rect 221 597 255 631
rect 289 597 323 631
rect 357 597 391 631
rect 425 597 459 631
rect 493 597 527 631
rect 561 597 595 631
rect 629 597 663 631
rect -778 493 -744 527
rect -778 425 -744 459
rect -778 357 -744 391
rect -778 289 -744 323
rect -778 221 -744 255
rect -778 153 -744 187
rect -778 85 -744 119
rect -778 17 -744 51
rect -778 -51 -744 -17
rect -778 -119 -744 -85
rect -778 -187 -744 -153
rect -778 -255 -744 -221
rect -778 -323 -744 -289
rect -778 -391 -744 -357
rect -778 -459 -744 -425
rect -778 -527 -744 -493
rect 744 493 778 527
rect 744 425 778 459
rect 744 357 778 391
rect 744 289 778 323
rect 744 221 778 255
rect 744 153 778 187
rect 744 85 778 119
rect 744 17 778 51
rect 744 -51 778 -17
rect 744 -119 778 -85
rect 744 -187 778 -153
rect 744 -255 778 -221
rect 744 -323 778 -289
rect 744 -391 778 -357
rect 744 -459 778 -425
rect 744 -527 778 -493
rect -663 -631 -629 -597
rect -595 -631 -561 -597
rect -527 -631 -493 -597
rect -459 -631 -425 -597
rect -391 -631 -357 -597
rect -323 -631 -289 -597
rect -255 -631 -221 -597
rect -187 -631 -153 -597
rect -119 -631 -85 -597
rect -51 -631 -17 -597
rect 17 -631 51 -597
rect 85 -631 119 -597
rect 153 -631 187 -597
rect 221 -631 255 -597
rect 289 -631 323 -597
rect 357 -631 391 -597
rect 425 -631 459 -597
rect 493 -631 527 -597
rect 561 -631 595 -597
rect 629 -631 663 -597
<< xpolycontact >>
rect -648 69 -510 501
rect -648 -501 -510 -69
rect -262 69 -124 501
rect -262 -501 -124 -69
rect 124 69 262 501
rect 124 -501 262 -69
rect 510 69 648 501
rect 510 -501 648 -69
<< ppolyres >>
rect -648 -69 -510 69
rect -262 -69 -124 69
rect 124 -69 262 69
rect 510 -69 648 69
<< locali >>
rect -778 597 -663 631
rect -629 597 -595 631
rect -561 597 -527 631
rect -493 597 -459 631
rect -425 597 -391 631
rect -357 597 -323 631
rect -289 597 -255 631
rect -221 597 -187 631
rect -153 597 -119 631
rect -85 597 -51 631
rect -17 597 17 631
rect 51 597 85 631
rect 119 597 153 631
rect 187 597 221 631
rect 255 597 289 631
rect 323 597 357 631
rect 391 597 425 631
rect 459 597 493 631
rect 527 597 561 631
rect 595 597 629 631
rect 663 597 778 631
rect -778 527 -744 597
rect 744 527 778 597
rect -778 459 -744 493
rect -778 391 -744 425
rect -778 323 -744 357
rect -778 255 -744 289
rect -778 187 -744 221
rect -778 119 -744 153
rect -778 51 -744 85
rect 744 459 778 493
rect 744 391 778 425
rect 744 323 778 357
rect 744 255 778 289
rect 744 187 778 221
rect 744 119 778 153
rect -778 -17 -744 17
rect -778 -85 -744 -51
rect 744 51 778 85
rect 744 -17 778 17
rect -778 -153 -744 -119
rect -778 -221 -744 -187
rect -778 -289 -744 -255
rect -778 -357 -744 -323
rect -778 -425 -744 -391
rect -778 -493 -744 -459
rect 744 -85 778 -51
rect 744 -153 778 -119
rect 744 -221 778 -187
rect 744 -289 778 -255
rect 744 -357 778 -323
rect 744 -425 778 -391
rect 744 -493 778 -459
rect -778 -597 -744 -527
rect 744 -597 778 -527
rect -778 -631 -663 -597
rect -629 -631 -595 -597
rect -561 -631 -527 -597
rect -493 -631 -459 -597
rect -425 -631 -391 -597
rect -357 -631 -323 -597
rect -289 -631 -255 -597
rect -221 -631 -187 -597
rect -153 -631 -119 -597
rect -85 -631 -51 -597
rect -17 -631 17 -597
rect 51 -631 85 -597
rect 119 -631 153 -597
rect 187 -631 221 -597
rect 255 -631 289 -597
rect 323 -631 357 -597
rect 391 -631 425 -597
rect 459 -631 493 -597
rect 527 -631 561 -597
rect 595 -631 629 -597
rect 663 -631 778 -597
<< viali >>
rect -632 87 -526 481
rect -246 87 -140 481
rect 140 87 246 481
rect 526 87 632 481
rect -632 -482 -526 -88
rect -246 -482 -140 -88
rect 140 -482 246 -88
rect 526 -482 632 -88
<< metal1 >>
rect -638 481 -520 495
rect -638 87 -632 481
rect -526 87 -520 481
rect -638 74 -520 87
rect -252 481 -134 495
rect -252 87 -246 481
rect -140 87 -134 481
rect -252 74 -134 87
rect 134 481 252 495
rect 134 87 140 481
rect 246 87 252 481
rect 134 74 252 87
rect 520 481 638 495
rect 520 87 526 481
rect 632 87 638 481
rect 520 74 638 87
rect -638 -88 -520 -74
rect -638 -482 -632 -88
rect -526 -482 -520 -88
rect -638 -495 -520 -482
rect -252 -88 -134 -74
rect -252 -482 -246 -88
rect -140 -482 -134 -88
rect -252 -495 -134 -482
rect 134 -88 252 -74
rect 134 -482 140 -88
rect 246 -482 252 -88
rect 134 -495 252 -482
rect 520 -88 638 -74
rect 520 -482 526 -88
rect 632 -482 638 -88
rect 520 -495 638 -482
<< properties >>
string FIXED_BBOX -761 -614 761 614
<< end >>
