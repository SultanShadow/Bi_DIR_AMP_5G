magic
tech sky130A
magscale 1 2
timestamp 1634927741
<< pwell >>
rect -191 1502 191 1588
rect -191 -1502 -105 1502
rect 105 -1502 191 1502
rect -191 -1588 191 -1502
<< psubdiff >>
rect -165 1528 -51 1562
rect -17 1528 17 1562
rect 51 1528 165 1562
rect -165 1445 -131 1528
rect 131 1445 165 1528
rect -165 1377 -131 1411
rect -165 1309 -131 1343
rect -165 1241 -131 1275
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect -165 -1275 -131 -1241
rect -165 -1343 -131 -1309
rect -165 -1411 -131 -1377
rect 131 1377 165 1411
rect 131 1309 165 1343
rect 131 1241 165 1275
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect 131 -1275 165 -1241
rect 131 -1343 165 -1309
rect 131 -1411 165 -1377
rect -165 -1528 -131 -1445
rect 131 -1528 165 -1445
rect -165 -1562 -51 -1528
rect -17 -1562 17 -1528
rect 51 -1562 165 -1528
<< psubdiffcont >>
rect -51 1528 -17 1562
rect 17 1528 51 1562
rect -165 1411 -131 1445
rect -165 1343 -131 1377
rect -165 1275 -131 1309
rect -165 1207 -131 1241
rect -165 1139 -131 1173
rect -165 1071 -131 1105
rect -165 1003 -131 1037
rect -165 935 -131 969
rect -165 867 -131 901
rect -165 799 -131 833
rect -165 731 -131 765
rect -165 663 -131 697
rect -165 595 -131 629
rect -165 527 -131 561
rect -165 459 -131 493
rect -165 391 -131 425
rect -165 323 -131 357
rect -165 255 -131 289
rect -165 187 -131 221
rect -165 119 -131 153
rect -165 51 -131 85
rect -165 -17 -131 17
rect -165 -85 -131 -51
rect -165 -153 -131 -119
rect -165 -221 -131 -187
rect -165 -289 -131 -255
rect -165 -357 -131 -323
rect -165 -425 -131 -391
rect -165 -493 -131 -459
rect -165 -561 -131 -527
rect -165 -629 -131 -595
rect -165 -697 -131 -663
rect -165 -765 -131 -731
rect -165 -833 -131 -799
rect -165 -901 -131 -867
rect -165 -969 -131 -935
rect -165 -1037 -131 -1003
rect -165 -1105 -131 -1071
rect -165 -1173 -131 -1139
rect -165 -1241 -131 -1207
rect -165 -1309 -131 -1275
rect -165 -1377 -131 -1343
rect -165 -1445 -131 -1411
rect 131 1411 165 1445
rect 131 1343 165 1377
rect 131 1275 165 1309
rect 131 1207 165 1241
rect 131 1139 165 1173
rect 131 1071 165 1105
rect 131 1003 165 1037
rect 131 935 165 969
rect 131 867 165 901
rect 131 799 165 833
rect 131 731 165 765
rect 131 663 165 697
rect 131 595 165 629
rect 131 527 165 561
rect 131 459 165 493
rect 131 391 165 425
rect 131 323 165 357
rect 131 255 165 289
rect 131 187 165 221
rect 131 119 165 153
rect 131 51 165 85
rect 131 -17 165 17
rect 131 -85 165 -51
rect 131 -153 165 -119
rect 131 -221 165 -187
rect 131 -289 165 -255
rect 131 -357 165 -323
rect 131 -425 165 -391
rect 131 -493 165 -459
rect 131 -561 165 -527
rect 131 -629 165 -595
rect 131 -697 165 -663
rect 131 -765 165 -731
rect 131 -833 165 -799
rect 131 -901 165 -867
rect 131 -969 165 -935
rect 131 -1037 165 -1003
rect 131 -1105 165 -1071
rect 131 -1173 165 -1139
rect 131 -1241 165 -1207
rect 131 -1309 165 -1275
rect 131 -1377 165 -1343
rect 131 -1445 165 -1411
rect -51 -1562 -17 -1528
rect 17 -1562 51 -1528
<< xpolycontact >>
rect -35 1000 35 1432
rect -35 -1432 35 -1000
<< ppolyres >>
rect -35 -1000 35 1000
<< locali >>
rect -165 1528 -51 1562
rect -17 1528 17 1562
rect 51 1528 165 1562
rect -165 1445 -131 1528
rect 131 1445 165 1528
rect -165 1377 -131 1411
rect -165 1309 -131 1343
rect -165 1241 -131 1275
rect -165 1173 -131 1207
rect -165 1105 -131 1139
rect -165 1037 -131 1071
rect -165 969 -131 1003
rect 131 1377 165 1411
rect 131 1309 165 1343
rect 131 1241 165 1275
rect 131 1173 165 1207
rect 131 1105 165 1139
rect 131 1037 165 1071
rect -165 901 -131 935
rect -165 833 -131 867
rect -165 765 -131 799
rect -165 697 -131 731
rect -165 629 -131 663
rect -165 561 -131 595
rect -165 493 -131 527
rect -165 425 -131 459
rect -165 357 -131 391
rect -165 289 -131 323
rect -165 221 -131 255
rect -165 153 -131 187
rect -165 85 -131 119
rect -165 17 -131 51
rect -165 -51 -131 -17
rect -165 -119 -131 -85
rect -165 -187 -131 -153
rect -165 -255 -131 -221
rect -165 -323 -131 -289
rect -165 -391 -131 -357
rect -165 -459 -131 -425
rect -165 -527 -131 -493
rect -165 -595 -131 -561
rect -165 -663 -131 -629
rect -165 -731 -131 -697
rect -165 -799 -131 -765
rect -165 -867 -131 -833
rect -165 -935 -131 -901
rect -165 -1003 -131 -969
rect 131 969 165 1003
rect 131 901 165 935
rect 131 833 165 867
rect 131 765 165 799
rect 131 697 165 731
rect 131 629 165 663
rect 131 561 165 595
rect 131 493 165 527
rect 131 425 165 459
rect 131 357 165 391
rect 131 289 165 323
rect 131 221 165 255
rect 131 153 165 187
rect 131 85 165 119
rect 131 17 165 51
rect 131 -51 165 -17
rect 131 -119 165 -85
rect 131 -187 165 -153
rect 131 -255 165 -221
rect 131 -323 165 -289
rect 131 -391 165 -357
rect 131 -459 165 -425
rect 131 -527 165 -493
rect 131 -595 165 -561
rect 131 -663 165 -629
rect 131 -731 165 -697
rect 131 -799 165 -765
rect 131 -867 165 -833
rect 131 -935 165 -901
rect -165 -1071 -131 -1037
rect -165 -1139 -131 -1105
rect -165 -1207 -131 -1173
rect -165 -1275 -131 -1241
rect -165 -1343 -131 -1309
rect -165 -1411 -131 -1377
rect 131 -1003 165 -969
rect 131 -1071 165 -1037
rect 131 -1139 165 -1105
rect 131 -1207 165 -1173
rect 131 -1275 165 -1241
rect 131 -1343 165 -1309
rect 131 -1411 165 -1377
rect -165 -1528 -131 -1445
rect 131 -1528 165 -1445
rect -165 -1562 -51 -1528
rect -17 -1562 17 -1528
rect 51 -1562 165 -1528
<< viali >>
rect -17 1378 17 1412
rect -17 1306 17 1340
rect -17 1234 17 1268
rect -17 1162 17 1196
rect -17 1090 17 1124
rect -17 1018 17 1052
rect -17 -1053 17 -1019
rect -17 -1125 17 -1091
rect -17 -1197 17 -1163
rect -17 -1269 17 -1235
rect -17 -1341 17 -1307
rect -17 -1413 17 -1379
<< metal1 >>
rect -25 1412 25 1426
rect -25 1378 -17 1412
rect 17 1378 25 1412
rect -25 1340 25 1378
rect -25 1306 -17 1340
rect 17 1306 25 1340
rect -25 1268 25 1306
rect -25 1234 -17 1268
rect 17 1234 25 1268
rect -25 1196 25 1234
rect -25 1162 -17 1196
rect 17 1162 25 1196
rect -25 1124 25 1162
rect -25 1090 -17 1124
rect 17 1090 25 1124
rect -25 1052 25 1090
rect -25 1018 -17 1052
rect 17 1018 25 1052
rect -25 1005 25 1018
rect -25 -1019 25 -1005
rect -25 -1053 -17 -1019
rect 17 -1053 25 -1019
rect -25 -1091 25 -1053
rect -25 -1125 -17 -1091
rect 17 -1125 25 -1091
rect -25 -1163 25 -1125
rect -25 -1197 -17 -1163
rect 17 -1197 25 -1163
rect -25 -1235 25 -1197
rect -25 -1269 -17 -1235
rect 17 -1269 25 -1235
rect -25 -1307 25 -1269
rect -25 -1341 -17 -1307
rect 17 -1341 25 -1307
rect -25 -1379 25 -1341
rect -25 -1413 -17 -1379
rect 17 -1413 25 -1379
rect -25 -1426 25 -1413
<< properties >>
string FIXED_BBOX -148 -1545 148 1545
<< end >>
