magic
tech sky130A
magscale 1 2
timestamp 1634906159
<< pwell >>
rect 9068 5733 9096 5740
<< locali >>
rect 6239 21889 6632 22186
rect 9068 21889 9341 21898
rect 6239 21886 9341 21889
rect 6240 20081 9341 21886
rect 9068 12151 9341 20081
rect 8251 10317 9292 10790
rect 8251 7547 9663 10317
rect 7675 -777 8880 278
rect 21710 147 21766 301
rect 22279 147 22336 301
rect 21710 113 22336 147
rect 7675 -953 7751 -777
rect 8808 -953 8880 -777
rect 7675 -1008 8880 -953
<< viali >>
rect 21766 147 22279 324
rect 7751 -953 8808 -777
<< metal1 >>
rect 10100 20801 10686 22109
rect 10100 20587 10230 20801
rect 10590 20587 10686 20801
rect 10100 20465 10686 20587
rect 20916 20803 22367 20923
rect 20916 20565 21183 20803
rect 22140 20565 22367 20803
rect 16137 19908 16203 19932
rect 20916 19807 22367 20565
rect 20916 19680 22363 19807
rect 20916 19255 21024 19680
rect 22241 19255 22363 19680
rect 4746 11413 4769 11548
rect 18350 11430 18372 11611
rect 20916 7963 22363 19255
rect 20916 7851 22626 7963
rect 20916 7250 21100 7851
rect 22198 7250 22626 7851
rect 20916 7115 22626 7250
rect 24154 7531 25284 7716
rect 24154 7088 24432 7531
rect 25084 7088 25284 7531
rect 25714 7231 26132 7265
rect 24154 6862 25284 7088
rect 9299 6447 25286 6862
rect 9068 5733 9096 5740
rect 6847 3355 6851 3373
rect 14495 1810 14806 4002
rect 11512 1551 11518 1617
rect 7796 1407 13978 1473
rect 7796 1058 13344 1407
rect 10586 385 10590 455
rect 13282 -236 13344 1058
rect 13903 -236 13978 1407
rect 17168 192 17605 391
rect 21669 324 22340 386
rect 13282 -292 13978 -236
rect 21669 147 21766 324
rect 22279 147 22340 324
rect 21669 -704 22340 147
rect 23385 45 23833 52
rect 23385 13 23833 29
rect 17168 -707 22340 -704
rect 7675 -777 22340 -707
rect 7675 -953 7751 -777
rect 8808 -953 22340 -777
rect 7675 -1008 22340 -953
<< via1 >>
rect 10230 20587 10590 20801
rect 21183 20565 22140 20803
rect 21024 19255 22241 19680
rect 21100 7250 22198 7851
rect 24432 7088 25084 7531
rect 13344 -236 13903 1407
<< metal2 >>
rect 3161 21130 3210 21778
rect 20783 20916 22367 20923
rect 6644 20803 22367 20916
rect 6644 20801 21183 20803
rect 6644 20587 10230 20801
rect 10590 20587 21183 20801
rect 6644 20565 21183 20587
rect 22140 20565 22367 20803
rect 6644 20465 22367 20565
rect 16989 20059 17135 20076
rect 18489 19680 22363 19808
rect 18489 19255 21024 19680
rect 22241 19255 22363 19680
rect 18489 19142 22363 19255
rect 9900 16872 11015 17236
rect 9900 13232 10206 16872
rect 10755 13232 11015 16872
rect 9900 12902 11015 13232
rect 11647 13328 18207 13554
rect 11647 12991 14236 13328
rect 17195 12991 18207 13328
rect 11647 12869 18207 12991
rect 10511 9670 19534 9763
rect 10511 9221 18109 9670
rect 18983 9221 19534 9670
rect 10511 9115 19534 9221
rect 11424 7851 22630 7965
rect 11424 7250 21100 7851
rect 22198 7250 22630 7851
rect 11424 7115 22630 7250
rect 23139 7667 23744 7784
rect 23139 7320 23269 7667
rect 23616 7320 23744 7667
rect 23139 6948 23744 7320
rect 24154 7531 25284 7716
rect 24154 7088 24432 7531
rect 25084 7088 25284 7531
rect 24154 7021 25284 7088
rect 17187 2947 18219 2955
rect 12450 1979 19290 2947
rect 17187 1529 18219 1979
rect 13282 1407 13978 1473
rect 13282 -236 13344 1407
rect 13903 -236 13978 1407
rect 13282 -292 13978 -236
<< via2 >>
rect 10206 13232 10755 16872
rect 14236 12991 17195 13328
rect 18109 9221 18983 9670
rect 23269 7320 23616 7667
rect 24432 7088 25084 7531
rect 13344 -236 13903 1407
<< metal3 >>
rect 9899 16872 11015 17237
rect 9899 13232 10206 16872
rect 10755 13232 11015 16872
rect 9899 12902 11015 13232
rect 13560 13328 18058 13554
rect 13560 12991 14236 13328
rect 17195 12991 18058 13328
rect 13560 12869 18058 12991
rect 18012 9670 19175 9763
rect 18012 9221 18109 9670
rect 18983 9221 19175 9670
rect 18012 9115 19175 9221
rect 23139 7667 23744 7784
rect 23139 7320 23269 7667
rect 23616 7320 23744 7667
rect 23139 7203 23744 7320
rect 24154 7531 25284 7716
rect 24154 7088 24432 7531
rect 25084 7088 25284 7531
rect 24154 7021 25284 7088
rect 13282 1407 13978 1473
rect 13282 -236 13344 1407
rect 13903 -236 13978 1407
rect 13282 -292 13978 -236
<< via3 >>
rect 10206 13232 10755 16872
rect 14236 12991 17195 13328
rect 18109 9221 18983 9670
rect 23269 7320 23616 7667
rect 24432 7088 25084 7531
rect 13344 -236 13903 1407
<< metal4 >>
rect 9899 16872 11015 17237
rect 9899 13232 10206 16872
rect 10755 13232 11015 16872
rect 9899 12902 11015 13232
rect 13560 13328 18058 13554
rect 13560 12991 14236 13328
rect 17195 12991 18058 13328
rect 13560 12869 18058 12991
rect 18012 9670 19576 9763
rect 18012 9221 18109 9670
rect 18983 9221 19576 9670
rect 18012 9115 19576 9221
rect 23139 7667 23744 7784
rect 23139 7320 23269 7667
rect 23616 7320 23744 7667
rect 23139 7203 23744 7320
rect 24154 7531 25284 7716
rect 24154 7088 24432 7531
rect 25084 7088 25284 7531
rect 24154 7021 25284 7088
rect 13282 1407 13978 1473
rect 13282 -236 13344 1407
rect 13903 -236 13978 1407
rect 13282 -292 13978 -236
<< via4 >>
rect 14236 12991 17195 13328
rect 23269 7320 23616 7667
rect 24432 7088 25084 7531
rect 13344 -236 13903 1407
<< metal5 >>
rect 13560 13328 18058 15016
rect 13560 12991 14236 13328
rect 17195 12991 18058 13328
rect 13560 12869 18058 12991
rect 18064 9115 19576 9763
rect 23139 7667 23744 8578
rect 23139 7320 23269 7667
rect 23616 7320 23744 7667
rect 23139 7203 23744 7320
rect 24154 7531 25284 7716
rect 24154 7088 24432 7531
rect 25084 7088 25284 7531
rect 24154 6650 25284 7088
rect 13282 1407 15152 1473
rect 13282 -236 13344 1407
rect 13903 -236 15152 1407
rect 13282 -292 15152 -236
use LNA  LNA_0
timestamp 1634905962
transform 1 0 6847 0 1 2730
box -6847 -2730 6094 5235
use LNA_Buff  LNA_Buff_0
timestamp 1634905962
transform -1 0 18309 0 1 18676
box -476 -5034 6978 1638
use sky130_fd_pr__cap_mim_m3_2_LJ5JLG  sky130_fd_pr__cap_mim_m3_2_LJ5JLG_0
timestamp 1634905962
transform -1 0 22629 0 1 11359
box -3351 -3101 3373 3101
use LNA_2ndstage  LNA_2ndstage_0
timestamp 1634905962
transform 1 0 20364 0 1 902
box -6280 -889 7501 7084
use Switch  Switch_0
timestamp 1634904720
transform 1 0 10953 0 1 9891
box -6207 -129 7419 3455
use PA_BUFF  PA_BUFF_0
timestamp 1634905962
transform 1 0 3802 0 -1 21092
box -641 -1250 6968 8136
<< labels >>
rlabel metal1 4747 11473 4747 11473 1 VSWN
rlabel metal1 18368 11505 18368 11505 1 VSWP
rlabel metal1 10685 21626 10685 21626 1 VDD
rlabel metal1 11517 1585 11517 1585 1 VBIAS1
rlabel metal1 9082 5739 9082 5739 1 VSS
rlabel metal1 6847 3362 6847 3362 1 VCASC1
rlabel metal1 10589 416 10589 416 1 VBIAS2
rlabel metal1 23636 16 23636 16 1 VBIAS3
rlabel metal1 25902 7253 25902 7253 1 VCASC2
rlabel metal2 17068 20074 17068 20074 1 RFOUTLNA
rlabel metal1 16171 19930 16171 19930 1 VBIAS4
rlabel metal2 3161 21423 3161 21423 1 RFOUTPA
<< end >>
